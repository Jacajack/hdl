`include "tb_common.svh"

module simple_dma_tb;
	initial begin
		`START_DUMP(simple_dma_tb);
	end
endmodule
